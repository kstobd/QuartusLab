module AndGate_Verilog (
    input A,
    input B,
    output Y
);
    assign Y = A & B;
endmodule
