VHDL code